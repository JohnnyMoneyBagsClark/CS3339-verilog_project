// nand_gate.v
module nand_gate (
    input wire [3:0] a,
    input wire [3:0] b,
    output wire [3:0] y
);
    assign y = ~(a & b);  // Vectorized NAND operation
endmodule

